///////////////////////////////////////////////////////////////////////////////
//   __  __          _____      _         _   _  ______      _______ _____   //
//  |  \/  |   /\   |  __ \    | |  /\   | \ | |/ __ \ \    / /_   _/ ____|  //
//  | \  / |  /  \  | |__) |   | | /  \  |  \| | |  | \ \  / /  | || |       //
//  | |\/| | / /\ \ |  _  /_   | |/ /\ \ | . ` | |  | |\ \/ /   | || |       //
//  | |  | |/ ____ \| | \ \ |__| / ____ \| |\  | |__| | \  /   _| || |____   //
//  |_|  |_/_/    \_\_|  \_\____/_/    \_\_| \_|\____/   \/   |_____\_____|  //
//                                                                           //
//                          JAN MARJANOVIC, 2014                             //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns/100ps

module cart_capture_tb;

bit		clk = 0;
bit		reset = 0;

wire	[15:0]	cart_ad;
wire			cart_rd;
wire			cart_alel;
wire			cart_aleh;

wire	[31:0] 	addr_o;
wire	[31:0]	data_o;
wire			valid_o;

//=============================================================================
always #20 clk = !clk;

initial begin
	#100;
	reset = 1;
	#100;
	reset = 0; 
end

//=============================================================================
cart_comm_wform cart_comm_wform_inst ( .* );

cart_capture cart_capture ( .* );

//=============================================================================
initial begin
	$display(" ---------------------------------------------- "); 
	$display("          Cartridge capture tesetbench          ");
	$display(" ---------------------------------------------- ");

	#(20us);
	$stop();
end


endmodule
