///////////////////////////////////////////////////////////////////////////////
//   __  __          _____      _         _   _  ______      _______ _____   //
//  |  \/  |   /\   |  __ \    | |  /\   | \ | |/ __ \ \    / /_   _/ ____|  //
//  | \  / |  /  \  | |__) |   | | /  \  |  \| | |  | \ \  / /  | || |       //
//  | |\/| | / /\ \ |  _  /_   | |/ /\ \ | . ` | |  | |\ \/ /   | || |       //
//  | |  | |/ ____ \| | \ \ |__| / ____ \| |\  | |__| | \  /   _| || |____   //
//  |_|  |_/_/    \_\_|  \_\____/_/    \_\_| \_|\____/   \/   |_____\_____|  //
//                                                                           //
//                          JAN MARJANOVIC, 2014                             //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns/100ps

module reset_gen # (
	parameter NR_CLK_CYCLES = 1_000_000
)(
	input		clk,	
	output reg		reset
);

reg [31:0] rst_cntr = 0;

always @ (posedge clk) begin
	if (rst_cntr < NR_CLK_CYCLES) begin
		rst_cntr	<= rst_cntr + 1;
		reset	<= 1'b1;
	end else begin
		reset	<= 1'b0;
	end
end

endmodule
